module jpeg_package();

endmodule 