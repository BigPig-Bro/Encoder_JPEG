module top(
    input           sys_clk,
    input           rst_n,

    input           start,

    // output          uart_tx

    output          send_data_vaild,send_data_last,
    output [7:0]    send_data
);

parameter   CLK_FRE         = 50_000_000; // sys_clk 时钟频率 50MHz\

parameter   H_ACTIVE        = 720; //编码图像宽度
parameter   V_ACTIVE        = 480; //编码图像高度


/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 		        测试输入源信号 	         /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
wire                rgb_clk, rgb_de;
wire [23:0]         rgb_data;

rgb_test #(
    .H_ACTIVE               (H_ACTIVE                   ),
    .V_ACTIVE               (V_ACTIVE                   )
)rgb_test_m0(
    .clk                    (sys_clk                    ),
    .rst_n                  (rst_n                      ),

    .start                  (start                      ),

    .rgb_clk                (rgb_clk                    ),
    .rgb_de                 (rgb_de                     ),
    .rgb_data               (rgb_data                   )
);

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			 Encoder_Jpeg 	            /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
// wire                send_data_vaild, send_data_last;
// wire [7:0]          send_data;

Encoder_Jpeg #(
    .H_ACTIVE               (H_ACTIVE                   ),
    .V_ACTIVE               (V_ACTIVE                   )
)Encoder_Jpeg_m0(
    .rst_n                  (rst_n                      ),
    .start                  (start                      ),

    .rgb_clk                (rgb_clk                    ),
    .rgb_de                 (rgb_de                     ),
    .rgb_data               (rgb_data                   ),

    .send_data_last         (send_data_last             ),
    .send_data_vaild        (send_data_vaild            ),
    .send_data              (send_data                  )
);

// /////////////////////////////////////////////////////////////////////////////////////////
// /////////////////////////////////////////////////////////////////////////////////////////
// //////////////////// 			  Uart 2 PC 	            /////////////////////////////
// /////////////////////////////////////////////////////////////////////////////////////////
// /////////////////////////////////////////////////////////////////////////////////////////
// uart_jpeg_top#(
//     .CLK_FRE                (CLK_FRE                    ),
//     .BAUD_RATE              (115200                     )
// )uart_jpeg_top_m0(
//     .clk                    (sys_clk                    ),

//     .send_data_vaild        (send_data_vaild            ),
//     .send_data              (send_data                  ),

//     .uart_tx                (uart_tx                    )
// );

endmodule 